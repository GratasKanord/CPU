module dmem (
    input  wire        clk,
    input  wire        rst,
    input  wire        we_dmem,          // Write enable (store)
    input  wire        is_LOAD,          // Load operation
    input  wire [7:0]  dmem_word_sel,    // Selects operation size
    input  wire [63:0] r_dmem_addr,      // Effective address
    input  wire [63:0] w_dmem_data,      // Data to write
    input  wire [2:0]  func3,            // Decoded command
    output reg  [63:0] dmem_data,        // Data to read
    output reg         exc_en,           // Exception enable
    output reg  [3:0]  exc_code,         // Exception code
    output reg  [63:0] exc_val           // Exception value (faulting address)
);

    localparam DMEM_SIZE = 16384;        // Increased to 16KB
    localparam DMEM_BASE = 64'h80000000; // Base address for memory mapping
    reg [7:0] dmem [0:DMEM_SIZE-1];      // Byte-addressable memory
    
    // Calculate offset address (subtract base to get local address)
    wire [63:0] local_addr = r_dmem_addr - DMEM_BASE;

    // Function to determine number of bytes per operation
    function integer get_num_bytes(input [7:0] sel);
        begin
            case (sel)
                8'b0000_0001: get_num_bytes = 1; // LB / SB
                8'b0000_0011: get_num_bytes = 2; // LH / SH
                8'b0000_1111: get_num_bytes = 4; // LW / SW
                8'b1111_1111: get_num_bytes = 8; // LD / SD
                default:      get_num_bytes = 1;
            endcase
        end
    endfunction

    // Memory initialization (for simulation)
    integer i, b;
    initial begin
        // Initialize all memory to zero first
        for (i = 0; i < DMEM_SIZE; i = i + 1)
            dmem[i] = 8'b0;
        
        // First, set the debug pattern
        for (i = 32'h2000; i < 32'h2020; i = i + 4) begin
            // Put address-dependent pattern
            dmem[i]   = i[7:0];      // LSB of address
            dmem[i+1] = i[15:8];     // Next byte
            dmem[i+2] = 8'hde;       // Debug pattern
            dmem[i+3] = 8'had;       // Debug pattern
        end
            
        dmem[32'h2006] = 8'hef;  
        dmem[32'h2007] = 8'hbe;  
            
        dmem[32'h2012] = 8'hef;
        dmem[32'h2013] = 8'hbe;
        dmem[32'h2014] = 8'h00;
        dmem[32'h2015] = 8'h00;

    end

    // Combinational: exception detection + load data output
    reg [3:0] num_bytes;

    always @(*) begin
        // Defaults
        exc_en   = 0;
        exc_code = 0;
        exc_val  = 0;
        dmem_data = 64'b0;

        num_bytes = get_num_bytes(dmem_word_sel);

        // Check if address is in our mapped range using local_addr
        if (r_dmem_addr < DMEM_BASE || local_addr >= DMEM_SIZE) begin
            if (we_dmem) begin
                exc_en   = 1;
                exc_code = 4'd7; // Store access fault
                exc_val  = r_dmem_addr;
            end else if (is_LOAD) begin
                exc_en   = 1;
                exc_code = 4'd5; // Load access fault  
                exc_val  = r_dmem_addr;
            end
        end
        // Check if the access would go beyond memory bounds
        else if (local_addr + num_bytes > DMEM_SIZE) begin
            if (we_dmem) begin
                exc_en   = 1;
                exc_code = 4'd7; // Store access fault
                exc_val  = r_dmem_addr;
            end else if (is_LOAD) begin
                exc_en   = 1;
                exc_code = 4'd5; // Load access fault  
                exc_val  = r_dmem_addr;
            end
        end
        // Check alignment (using original address for alignment checks)
        else if ((num_bytes == 2 && r_dmem_addr[0] != 0) ||
                 (num_bytes == 4 && r_dmem_addr[1:0] != 0) ||
                 (num_bytes == 8 && r_dmem_addr[2:0] != 0)) begin
            if (we_dmem) begin
                exc_en   = 1;
                exc_code = 4'd6; // Store address misaligned
                exc_val  = r_dmem_addr;
            end else if (is_LOAD) begin
                exc_en   = 1;
                exc_code = 4'd4; // Load address misaligned
                exc_val  = r_dmem_addr;
            end
        end
        // Handle tohost writes (compliance test exit condition)
        else if (we_dmem && r_dmem_addr == 64'h80001000) begin
            $display("TEST COMPLETE, to_host was written!");
            $finish;
        end
        // Normal load operation
        else if (is_LOAD && !we_dmem) begin
            dmem_data = 0;
            for (b = 0; b < num_bytes; b = b + 1)
                dmem_data[b*8 +: 8] = dmem[local_addr + b];
            
            // Extension based on instruction type
            case (dmem_word_sel)
                8'b0000_0001: begin // Byte loads
                    case (func3)
                        3'b000: dmem_data = {{56{dmem_data[7]}}, dmem_data[7:0]}; // LB - sign extend
                        3'b100: dmem_data = {56'b0, dmem_data[7:0]};              // LBU - zero extend
                        default: dmem_data = {{56{dmem_data[7]}}, dmem_data[7:0]}; // default to signed
                    endcase
                end
                8'b0000_0011: begin // Halfword loads  
                    case (func3)
                        3'b001: dmem_data = {{48{dmem_data[15]}}, dmem_data[15:0]}; // LH - sign extend
                        3'b101: dmem_data = {48'b0, dmem_data[15:0]};               // LHU - zero extend
                        default: dmem_data = {{48{dmem_data[15]}}, dmem_data[15:0]}; // default to signed
                    endcase
                end
                8'b0000_1111: begin // Word loads
                    case (func3)
                        3'b010: dmem_data = {{32{dmem_data[31]}}, dmem_data[31:0]}; // LW - sign extend
                        3'b110: dmem_data = {32'b0, dmem_data[31:0]};               // LWU - zero extend
                        default: dmem_data = {{32{dmem_data[31]}}, dmem_data[31:0]}; // default to signed
                    endcase
                end
            endcase
        end
    end

    // Sequential: perform store only if no exception
    always @(posedge clk) begin
        if (we_dmem && !exc_en && r_dmem_addr != 64'h80001000) begin
            for (b = 0; b < num_bytes; b = b + 1)
                dmem[local_addr + b] <= w_dmem_data[b*8 +: 8];
        end
    end

endmodule